module adder (
    input wire [3:0] a, b,
    output wire [4:0] sum
);
    assign sum = a + b;
endmodule

